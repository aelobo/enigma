/**
 * library.vh
 *
 * Enigma Machine
 *
 * ECE 18-500
 * Carnegie Mellon University
 *
 * This is the library of standard components used by the enigma machine,
 * which includes both synchronous and combinational components.
 **/


/*----------------------------------------------------------------------------*
 *  Combinational Components                                                  *
 *----------------------------------------------------------------------------*/


/*----------------------------------------------------------------------------*
 *  Synchronous Components                                                    *
 *----------------------------------------------------------------------------*/