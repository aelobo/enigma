/**
 * internal_defines.vh
 *
 * Enigma Machine
 *
 * ECE 18-500
 * Carnegie Mellon University
 *
 * This contains the definitions of constants and types that are used by the
 * enigma machine, such as ...
**/

`ifndef INTERNAL_DEFINES_VH_
`define INTERNAL_DEFINES_VH_

/*----------------------------------------------------------------------------*
 *  Enumerated Types                                                          *
 *----------------------------------------------------------------------------*/
 